`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company       : Self-made
// Engineer      : Muhammad Abdur-Rehman Siddiqui
//
// Create Date   : 15:54:41 12/06/2020
// Design Name   :
// Module Name   : tb_ALU_microprocessor
// Project Name  : Single cycle 16-bit ARM Microprocessor
// Target Devices:
// Tool versions : ISE Design Suite 14.7
// Description   : Test bench for ALU module for the processor
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module tb_ALU_microprocessor;

// Inputs
reg alu_clk;
reg [ 5:0] alu_ctrl   ;
reg [31:0] in_1       ;
reg [31:0] in_2       ;

// Outputs
wire [31:0] alu_rslt  ;
wire [ 4:0] alu_checks;

// Instantiate the Unit Under Test (UUT)
ALU_microprocessor alu_mp_design (
  .alu_ctrl  (alu_ctrl  ), 
  .in_1      (in_1      ), 
  .in_2      (in_2      ), 
  .alu_clk   (alu_clk   ), 
  .alu_rslt  (alu_rslt  ), 
  .alu_checks(alu_checks)
);

// ALU module operates on a whopping 8.93 GHz clock frequency accurately generated by point precision
always #0.055555556 alu_clk = ~alu_clk;
  
initial begin
// Initialize Inputs
  alu_ctrl    = 0;
  in_1        = 0;
  in_2        = 0;
  alu_clk     = 0;

  // Stalling some 100 cycles
  repeat(100)@(posedge alu_clk);

  //Initial assignments for inputs
  @(posedge alu_clk);
  in_1        = 32'b0;
  in_2        = 32'b0;
  alu_ctrl    =  6'hx;
  
  //Maximum Input randomization
  repeat(10000)@(posedge alu_clk) begin
    in_1     = $urandom;
    in_2     = $urandom;
    alu_ctrl = $urandom;
    @(posedge alu_clk);
  end //repeat
end //initial
      
endmodule

